/* Procedurally generated decoder. 
 * Generated using decoderGen script.
 */
module Decoder_5_32(decode_in, decode_out);
	input[4:0] decode_in;
	output[31:0] decode_out;
	assign decode_out =
		decode_in == 0 ? 32'b00000000000000000000000000000001 :
		decode_in == 1 ? 32'b00000000000000000000000000000010 :
		decode_in == 2 ? 32'b00000000000000000000000000000100 :
		decode_in == 3 ? 32'b00000000000000000000000000001000 :
		decode_in == 4 ? 32'b00000000000000000000000000010000 :
		decode_in == 5 ? 32'b00000000000000000000000000100000 :
		decode_in == 6 ? 32'b00000000000000000000000001000000 :
		decode_in == 7 ? 32'b00000000000000000000000010000000 :
		decode_in == 8 ? 32'b00000000000000000000000100000000 :
		decode_in == 9 ? 32'b00000000000000000000001000000000 :
		decode_in == 10 ? 32'b00000000000000000000010000000000 :
		decode_in == 11 ? 32'b00000000000000000000100000000000 :
		decode_in == 12 ? 32'b00000000000000000001000000000000 :
		decode_in == 13 ? 32'b00000000000000000010000000000000 :
		decode_in == 14 ? 32'b00000000000000000100000000000000 :
		decode_in == 15 ? 32'b00000000000000001000000000000000 :
		decode_in == 16 ? 32'b00000000000000010000000000000000 :
		decode_in == 17 ? 32'b00000000000000100000000000000000 :
		decode_in == 18 ? 32'b00000000000001000000000000000000 :
		decode_in == 19 ? 32'b00000000000010000000000000000000 :
		decode_in == 20 ? 32'b00000000000100000000000000000000 :
		decode_in == 21 ? 32'b00000000001000000000000000000000 :
		decode_in == 22 ? 32'b00000000010000000000000000000000 :
		decode_in == 23 ? 32'b00000000100000000000000000000000 :
		decode_in == 24 ? 32'b00000001000000000000000000000000 :
		decode_in == 25 ? 32'b00000010000000000000000000000000 :
		decode_in == 26 ? 32'b00000100000000000000000000000000 :
		decode_in == 27 ? 32'b00001000000000000000000000000000 :
		decode_in == 28 ? 32'b00010000000000000000000000000000 :
		decode_in == 29 ? 32'b00100000000000000000000000000000 :
		decode_in == 30 ? 32'b01000000000000000000000000000000 :
		decode_in == 31 ? 32'b10000000000000000000000000000000 :
		0;
endmodule